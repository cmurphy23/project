module FreqLUT(input [7:0] message, output[9:0] freq);


   
endmodule
