`ifndef MIDI_MESSAGE
`define MIDI_MESSAGE

`define MIDI_NOTE_ON 4'b1001
`define MIDI_NOTE_OFF 4'b1000
`define MIDI_PITCH_WHEEL 4'b1110


`define MIDI_EVENT 2'b00
`define MIDI_FREQ 2'b01
`define MIDI_VEL 2'b10

`endif //MIDI_MESSAGE
